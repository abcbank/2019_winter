module Interpol(data_in_re, data_in_im, data_out_re, data_out_re);

input signed 